CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 30 400 10
176 80 1918 940
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
47 C:\Users\User\Desktop\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
17
4 LED~
171 328 122 0 2 2
10 6 2
0
0 0 864 0
4 LED0
22 22 50 30
1 S
28 -10 35 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
6421 0 0
2
44773.8 0
0
8 3-In OR~
219 270 111 0 4 22
0 5 7 4 6
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
7743 0 0
2
44773.8 0
0
9 Inverter~
13 140 171 0 2 22
0 8 9
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
9840 0 0
2
44773.8 0
0
9 Inverter~
13 143 50 0 2 22
0 8 11
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
6910 0 0
2
44773.8 0
0
9 Inverter~
13 146 88 0 2 22
0 8 3
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
449 0 0
2
44773.8 0
0
5 7415~
219 198 152 0 4 22
0 8 11 9 4
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 1 0
1 U
8761 0 0
2
44773.8 0
0
5 7415~
219 198 111 0 4 22
0 8 3 9 7
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
6748 0 0
2
44773.8 0
0
5 7415~
219 198 70 0 4 22
0 11 8 3 5
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 1 0
1 U
7393 0 0
2
44773.8 0
0
7 Ground~
168 328 139 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7699 0 0
2
44773.7 0
0
7 Ground~
168 87 81 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6638 0 0
2
44773.7 1
0
12 SPDT Switch~
164 104 70 0 10 11
0 8 8 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 A
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
4595 0 0
2
44773.7 0
0
7 Ground~
168 87 154 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9395 0 0
2
44773.7 1
0
12 SPDT Switch~
164 104 143 0 10 11
0 8 8 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 C
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3303 0 0
2
44773.7 0
0
7 Ground~
168 13 72 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4498 0 0
2
5.90041e-315 0
0
9 V Source~
197 45 65 0 2 5
0 8 2
0
0 0 17264 270
2 5V
-7 -20 7 -12
3 Vs1
-11 -30 10 -22
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
9728 0 0
2
5.90041e-315 0
0
7 Ground~
168 85 118 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3789 0 0
2
5.90041e-315 0
0
12 SPDT Switch~
164 102 107 0 10 11
0 8 8 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 B
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3978 0 0
2
5.90041e-315 0
0
24
2 0 3 0 0 4224 0 7 0 0 14 2
174 111
174 88
3 4 4 0 0 4224 0 2 6 0 0 3
257 120
219 120
219 152
1 4 5 0 0 4224 0 2 8 0 0 3
257 102
219 102
219 70
1 4 6 0 0 8320 0 1 2 0 0 3
328 112
328 111
303 111
2 4 7 0 0 4224 0 2 7 0 0 4
258 111
218 111
218 111
219 111
0 1 8 0 0 4096 0 0 7 12 0 2
119 102
174 102
3 2 9 0 0 8320 0 7 3 0 0 3
174 120
161 120
161 171
0 1 8 0 0 4224 10 0 3 15 0 2
125 70
125 171
0 2 11 0 0 4224 0 0 6 13 0 3
165 50
165 152
174 152
2 3 9 0 0 0 0 3 6 0 0 3
161 171
174 171
174 161
1 0 8 0 0 4224 12 5 0 0 16 2
131 88
131 143
1 1 8 0 0 8320 0 4 17 0 0 3
128 50
119 50
119 107
2 1 11 0 0 128 0 4 8 0 0 3
164 50
174 50
174 61
2 3 3 0 0 128 0 5 8 0 0 3
167 88
174 88
174 79
2 1 8 0 0 128 10 8 11 0 0 2
174 70
121 70
1 1 8 0 0 128 12 6 13 0 0 2
174 143
121 143
0 1 8 0 0 12288 13 0 15 20 0 4
66 103
66 101
65 101
65 66
1 2 2 0 0 4096 0 9 1 0 0 2
328 133
328 132
2 0 8 0 0 0 13 11 0 0 17 2
87 66
65 66
2 2 8 0 0 8320 13 17 13 0 0 4
85 103
65 103
65 139
87 139
2 1 2 0 0 4224 0 15 14 0 0 2
23 66
13 66
1 3 2 0 0 0 0 10 11 0 0 2
87 75
87 74
1 3 2 0 0 0 0 12 13 0 0 2
87 148
87 147
1 3 2 0 0 0 0 16 17 0 0 2
85 112
85 111
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
