CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 400 10
176 80 1918 940
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
47 C:\Users\User\Desktop\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
15
9 2-In XOR~
219 279 97 0 3 22
0 7 5 6
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
4797 0 0
2
44774.4 0
0
9 2-In XOR~
219 209 88 0 3 22
0 8 5 7
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4681 0 0
2
44774.4 0
0
9 2-In XOR~
219 149 79 0 3 22
0 5 5 8
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9730 0 0
2
44774.4 0
0
7 Ground~
168 87 187 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9874 0 0
2
44774.4 1
0
12 SPDT Switch~
164 104 176 0 10 11
0 5 5 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 D
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
364 0 0
2
44774.4 0
0
7 Ground~
168 86 152 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3656 0 0
2
44774.4 1
0
12 SPDT Switch~
164 103 141 0 10 11
0 5 5 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 C
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3131 0 0
2
44774.4 0
0
4 LED~
171 328 122 0 2 2
13 6 2
0
0 0 864 0
4 LED0
22 22 50 30
1 P
28 -10 35 -2
0
0
11 %D %1 %2 %M
0
0
0
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
6772 0 0
2
5.90041e-315 0
0
7 Ground~
168 328 139 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9557 0 0
2
5.90041e-315 0
0
7 Ground~
168 87 81 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5789 0 0
2
5.90041e-315 5.26354e-315
0
12 SPDT Switch~
164 104 70 0 10 11
0 5 5 2 0 0 0 0 0 0
1
0
0 0 4720 0
1 A
-4 -15 3 -7
1 A
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 -1 0
1 S
7328 0 0
2
5.90041e-315 0
0
7 Ground~
168 13 72 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4799 0 0
2
44773.8 0
0
9 V Source~
197 45 65 0 2 5
0 5 2
0
0 0 17264 270
2 5V
-7 -20 7 -12
3 Vs1
-11 -30 10 -22
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
9196 0 0
2
44773.8 1
0
7 Ground~
168 85 118 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3857 0 0
2
44773.8 2
0
12 SPDT Switch~
164 102 107 0 10 11
0 5 5 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 B
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
7125 0 0
2
44773.8 3
0
17
2 1 5 0 0 12416 3 1 5 0 0 4
263 106
241 106
241 176
121 176
2 1 5 0 0 12416 4 2 7 0 0 4
193 97
179 97
179 141
120 141
2 1 5 0 0 8320 0 3 15 0 0 3
133 88
119 88
119 107
3 1 6 0 0 4224 0 1 8 0 0 3
312 97
328 97
328 112
1 3 7 0 0 4224 0 1 2 0 0 2
263 88
242 88
1 3 8 0 0 4224 0 2 3 0 0 2
193 79
182 79
1 1 5 0 0 4224 9 3 11 0 0 2
133 70
121 70
2 0 5 0 0 8192 10 5 0 0 9 3
87 172
66 172
66 137
2 0 5 0 0 0 10 7 0 0 13 3
86 137
66 137
66 103
1 3 2 0 0 4096 0 4 5 0 0 2
87 181
87 180
1 3 2 0 0 0 0 6 7 0 0 2
86 146
86 145
2 1 5 0 0 0 10 11 13 0 0 2
87 66
65 66
2 1 5 0 0 8320 10 15 13 0 0 3
85 103
65 103
65 66
1 2 2 0 0 0 0 9 8 0 0 2
328 133
328 132
2 1 2 0 0 4224 0 13 12 0 0 2
23 66
13 66
1 3 2 0 0 0 0 10 11 0 0 2
87 75
87 74
1 3 2 0 0 0 0 14 15 0 0 2
85 112
85 111
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
