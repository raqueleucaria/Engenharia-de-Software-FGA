CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 400 10
176 80 1918 940
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
47 C:\Users\User\Desktop\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
18
9 Inverter~
13 136 143 0 2 22
0 6 4
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
5130 0 0
2
44773.8 0
0
9 Inverter~
13 186 104 0 2 22
0 5 7
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
391 0 0
2
44773.8 0
0
8 2-In OR~
219 285 62 0 3 22
0 11 9 10
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3124 0 0
2
44773.8 0
0
9 2-In AND~
219 230 138 0 3 22
0 5 4 3
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3421 0 0
2
44773.8 0
0
9 2-In AND~
219 230 95 0 3 22
0 6 7 9
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8157 0 0
2
44773.8 0
0
9 3-In AND~
219 230 53 0 4 22
0 6 5 4 11
0
0 0 624 0
5 74F11
-18 -28 17 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 1 0
1 U
5572 0 0
2
44773.8 0
0
7 Ground~
168 328 93 0 1 3
0 6
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8901 0 0
2
44773.8 1
0
4 LED~
171 328 76 0 2 2
10 10 6
0
0 0 864 0
4 LED0
22 22 50 30
2 B1
25 -10 39 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7361 0 0
2
44773.8 0
0
4 LED~
171 328 122 0 2 2
10 3 6
0
0 0 864 0
4 LED0
22 22 50 30
2 B2
25 -10 39 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4747 0 0
2
5.90041e-315 0
0
7 Ground~
168 328 139 0 1 3
0 6
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
972 0 0
2
5.90041e-315 0
0
7 Ground~
168 87 81 0 1 3
0 6
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3472 0 0
2
5.90041e-315 5.26354e-315
0
12 SPDT Switch~
164 104 70 0 3 11
0 6 5 6
0
0 0 4720 0
0
2 T1
-7 -16 7 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9998 0 0
2
5.90041e-315 0
0
7 Ground~
168 87 154 0 1 3
0 6
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3536 0 0
2
5.90041e-315 5.26354e-315
0
12 SPDT Switch~
164 104 143 0 3 11
0 6 5 6
0
0 0 4720 0
0
2 T3
-7 -16 7 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
4597 0 0
2
5.90041e-315 0
0
7 Ground~
168 13 72 0 1 3
0 6
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3835 0 0
2
44773.8 0
0
9 V Source~
197 45 65 0 2 5
0 5 6
0
0 0 17264 270
2 5V
-7 -20 7 -12
3 Vs1
-11 -30 10 -22
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
3670 0 0
2
44773.8 1
0
7 Ground~
168 85 118 0 1 3
0 6
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5616 0 0
2
44773.8 2
0
12 SPDT Switch~
164 102 107 0 10 11
0 5 5 6 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 T2
-7 -16 7 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9323 0 0
2
44773.8 3
0
22
1 3 3 0 0 4224 0 9 4 0 0 4
328 112
264 112
264 138
251 138
2 2 4 0 0 4096 0 4 1 0 0 3
206 147
157 147
157 143
1 0 5 0 0 4224 0 4 0 0 4 3
206 129
149 129
149 104
1 0 5 0 0 0 0 2 0 0 8 2
171 104
149 104
3 2 4 0 0 8320 0 6 1 0 0 3
206 62
157 62
157 143
1 1 6 0 0 0 0 1 14 0 0 2
121 143
121 143
2 2 7 0 0 4224 0 2 5 0 0 2
207 104
206 104
2 1 5 0 0 0 0 6 18 0 0 4
206 53
149 53
149 107
119 107
1 0 6 0 0 4224 8 5 0 0 10 3
206 86
138 86
138 70
1 1 6 0 0 0 8 12 6 0 0 4
121 70
138 70
138 44
206 44
2 3 9 0 0 8320 0 3 5 0 0 3
272 71
251 71
251 95
3 1 10 0 0 4224 0 3 8 0 0 3
318 62
328 62
328 66
1 4 11 0 0 4224 0 3 6 0 0 2
272 53
251 53
1 2 6 0 0 4112 2 7 8 0 0 2
328 87
328 86
0 1 5 0 0 12288 12 0 16 18 0 4
66 103
66 101
65 101
65 66
1 2 6 0 0 0 2 10 9 0 0 2
328 133
328 132
2 0 5 0 0 0 12 12 0 0 15 2
87 66
65 66
2 2 5 0 0 8320 12 18 14 0 0 4
85 103
65 103
65 139
87 139
2 1 6 0 0 4224 2 16 15 0 0 2
23 66
13 66
1 3 6 0 0 0 2 11 12 0 0 2
87 75
87 74
1 3 6 0 0 0 2 13 14 0 0 2
87 148
87 147
1 3 6 0 0 0 2 17 18 0 0 2
85 112
85 111
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
