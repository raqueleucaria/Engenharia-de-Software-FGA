CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 90 30 400 10
176 80 1918 940
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
47 C:\Users\User\Desktop\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
18
7 Ground~
168 32 188 0 1 3
0 9
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5130 0 0
2
44773.6 0
0
9 V Source~
197 32 162 0 2 5
0 3 9
0
0 0 17264 0
2 5V
16 0 30 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
391 0 0
2
44773.6 0
0
7 Ground~
168 235 134 0 1 3
0 9
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3124 0 0
2
44773.6 0
0
7 Ground~
168 234 176 0 1 3
0 9
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3421 0 0
2
44773.6 0
0
7 Ground~
168 234 221 0 1 3
0 9
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8157 0 0
2
44773.6 0
0
7 Ground~
168 84 227 0 1 3
0 9
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5572 0 0
2
44773.6 0
0
7 Ground~
168 84 175 0 1 3
0 9
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8901 0 0
2
44773.6 0
0
7 Ground~
168 85 118 0 1 3
0 9
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7361 0 0
2
44773.6 0
0
9 2-In AND~
219 199 196 0 3 22
0 6 5 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4747 0 0
2
44773.6 0
0
5 4049~
219 141 187 0 2 22
0 9 6
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
972 0 0
2
44773.6 0
0
5 4049~
219 141 141 0 2 22
0 9 5
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
3472 0 0
2
44773.6 0
0
12 SPDT Switch~
164 101 217 0 3 11
0 10 3 9
0
0 0 4720 0
0
1 C
-4 -15 3 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 512 0 0 0 0
1 S
9998 0 0
2
44773.6 0
0
12 SPDT Switch~
164 101 165 0 3 11
0 9 3 9
0
0 0 4720 0
0
1 B
-4 -15 3 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3536 0 0
2
44773.6 0
0
12 SPDT Switch~
164 102 108 0 3 11
0 9 3 9
0
0 0 4720 0
0
1 A
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
4597 0 0
2
44773.6 0
0
4 LED~
171 235 118 0 2 2
10 9 9
0
0 0 864 0
3 S_A
16 0 37 8
2 D3
20 -10 34 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3835 0 0
2
44773.6 0
0
4 LED~
171 234 160 0 2 2
10 8 9
0
0 0 864 0
3 S_B
20 0 41 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3670 0 0
2
44773.6 0
0
4 LED~
171 234 206 0 2 2
10 4 9
0
0 0 864 0
3 S_C
20 0 41 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
5616 0 0
2
44773.6 0
0
9 2-In AND~
219 198 150 0 3 22
0 5 9 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9323 0 0
2
44773.6 0
0
19
2 0 3 0 0 8192 0 12 0 0 2 3
84 213
67 213
67 161
2 0 3 0 0 0 0 13 0 0 3 4
84 161
67 161
67 135
32 135
2 1 3 0 0 4224 0 14 2 0 0 3
85 104
32 104
32 141
1 2 9 0 0 4224 2 1 2 0 0 2
32 182
32 183
1 2 9 0 0 0 2 3 15 0 0 2
235 128
235 128
1 2 9 0 0 0 2 4 16 0 0 2
234 170
234 170
1 2 9 0 0 128 2 5 17 0 0 2
234 215
234 216
1 3 9 0 0 0 2 6 12 0 0 2
84 221
84 221
1 3 9 0 0 0 2 7 13 0 0 2
84 169
84 169
1 3 9 0 0 0 2 8 14 0 0 2
85 112
85 112
3 1 4 0 0 4224 0 9 17 0 0 2
220 196
234 196
2 2 5 0 0 4224 0 11 9 0 0 3
162 141
162 205
175 205
2 1 6 0 0 4224 0 10 9 0 0 2
162 187
175 187
1 0 9 0 0 8192 7 10 0 0 18 3
126 187
121 187
121 165
3 1 8 0 0 4224 0 18 16 0 0 2
219 150
234 150
1 1 9 0 0 8192 0 11 14 0 0 3
126 141
119 141
119 108
2 1 5 0 0 0 0 11 18 0 0 2
162 141
174 141
1 2 9 0 0 4224 7 13 18 0 0 4
118 165
167 165
167 159
174 159
1 1 9 0 0 4224 0 14 15 0 0 2
119 108
235 108
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
