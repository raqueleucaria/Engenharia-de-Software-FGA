CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 60 30 400 10
176 80 1918 940
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
47 C:\Users\User\Desktop\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
9
7 Ground~
168 32 188 0 1 3
0 5
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
317 0 0
2
5.90041e-315 0
0
9 V Source~
197 32 162 0 2 5
0 4 5
0
0 0 17264 0
2 5V
16 0 30 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
3108 0 0
2
5.90041e-315 0
0
7 Ground~
168 235 134 0 1 3
0 5
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4299 0 0
2
5.90041e-315 0
0
7 Ground~
168 234 176 0 1 3
0 5
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9672 0 0
2
5.90041e-315 0
0
7 Ground~
168 85 118 0 1 3
0 5
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7876 0 0
2
5.90041e-315 0
0
5 4049~
219 141 141 0 2 22
0 5 3
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
6369 0 0
2
5.90041e-315 0
0
12 SPDT Switch~
164 102 107 0 3 11
0 5 4 5
0
0 0 4720 0
0
2 CA
-7 -16 7 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9172 0 0
2
5.90041e-315 0
0
4 LED~
171 235 117 0 2 2
10 5 5
0
0 0 880 0
3 S_A
16 0 37 8
2 D3
20 -10 34 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7100 0 0
2
5.90041e-315 0
0
4 LED~
171 234 160 0 2 2
10 3 5
0
0 0 880 0
3 S_B
20 0 41 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3820 0 0
2
5.90041e-315 0
0
8
2 1 3 0 0 4224 0 6 9 0 0 4
162 141
213 141
213 150
234 150
2 1 4 0 0 4224 0 7 2 0 0 3
85 103
32 103
32 141
1 2 5 0 0 4224 2 1 2 0 0 2
32 182
32 183
1 2 5 0 0 0 2 3 8 0 0 2
235 128
235 127
1 2 5 0 0 0 2 4 9 0 0 2
234 170
234 170
1 3 5 0 0 0 2 5 7 0 0 2
85 112
85 111
1 1 5 0 0 8192 0 6 7 0 0 3
126 141
119 141
119 107
1 1 5 0 0 4224 0 7 8 0 0 2
119 107
235 107
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
