CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 400 10
176 80 1918 940
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
47 C:\Users\User\Desktop\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
19
9 3-In AND~
219 265 134 0 4 22
0 4 4 5 8
0
0 0 624 0
5 74F11
-18 -28 17 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 4 0
1 U
7376 0 0
2
44774.4 0
0
8 2-In OR~
219 169 167 0 3 22
0 4 4 5
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9156 0 0
2
44774.4 0
0
9 Inverter~
13 207 84 0 2 22
0 4 9
0
0 0 112 0
5 74F04
-18 -19 17 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
5776 0 0
2
44774.4 0
0
9 Inverter~
13 207 48 0 2 22
0 4 10
0
0 0 112 0
5 74F04
-18 -19 17 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
7207 0 0
2
44774.4 0
0
9 2-In AND~
219 252 66 0 3 22
0 10 9 11
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4459 0 0
2
44774.4 0
0
7 Ground~
168 87 187 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3760 0 0
2
44774.4 1
0
12 SPDT Switch~
164 104 176 0 10 11
0 4 4 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 C
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
754 0 0
2
44774.4 0
0
7 Ground~
168 86 152 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9767 0 0
2
44774.4 1
0
12 SPDT Switch~
164 103 141 0 10 11
0 4 4 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 B
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
7978 0 0
2
44774.4 0
0
7 Ground~
168 328 93 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3142 0 0
2
44773.8 1
0
4 LED~
171 328 76 0 2 2
10 11 2
0
0 0 864 0
4 LED0
22 22 50 30
1 R
28 -10 35 -2
0
0
11 %D %1 %2 %M
0
0
0
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
3284 0 0
2
44773.8 0
0
4 LED~
171 328 122 0 2 2
12 8 2
0
0 0 864 0
4 LED0
22 22 50 30
1 G
28 -10 35 -2
0
0
11 %D %1 %2 %M
0
0
0
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
659 0 0
2
5.90041e-315 0
0
7 Ground~
168 328 139 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3800 0 0
2
5.90041e-315 0
0
7 Ground~
168 87 81 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6792 0 0
2
5.90041e-315 5.26354e-315
0
12 SPDT Switch~
164 104 70 0 10 11
0 4 4 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
4 MODO
-14 -16 14 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3701 0 0
2
5.90041e-315 0
0
7 Ground~
168 13 72 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6316 0 0
2
44773.8 0
0
9 V Source~
197 45 65 0 2 5
0 4 2
0
0 0 17264 270
2 5V
-7 -20 7 -12
3 Vs1
-11 -30 10 -22
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
8734 0 0
2
44773.8 1
0
7 Ground~
168 85 118 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7988 0 0
2
44773.8 2
0
12 SPDT Switch~
164 102 107 0 10 11
0 4 4 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 A
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3217 0 0
2
44773.8 3
0
22
0 1 4 0 0 8320 3 0 1 8 0 3
173 69
173 125
241 125
2 0 4 0 0 4224 0 1 0 0 7 3
241 134
150 134
150 107
3 3 5 0 0 4224 0 1 2 0 0 3
241 143
202 143
202 167
2 1 4 0 0 12416 6 2 7 0 0 4
156 176
157 176
157 176
121 176
1 1 4 0 0 4240 7 9 2 0 0 4
120 141
143 141
143 158
156 158
1 4 8 0 0 4224 0 12 1 0 0 3
328 112
286 112
286 134
1 1 4 0 0 0 0 3 19 0 0 4
192 84
150 84
150 107
119 107
1 1 4 0 0 0 3 4 15 0 0 4
192 48
173 48
173 70
121 70
2 2 9 0 0 4224 0 3 5 0 0 2
228 84
228 75
2 1 10 0 0 4224 0 4 5 0 0 2
228 48
228 57
3 1 11 0 0 4224 0 5 11 0 0 2
273 66
328 66
2 0 4 0 0 8192 12 7 0 0 13 3
87 172
66 172
66 137
2 0 4 0 0 0 12 9 0 0 17 3
86 137
66 137
66 103
1 3 2 0 0 4096 0 6 7 0 0 2
87 181
87 180
1 3 2 0 0 0 0 8 9 0 0 2
86 146
86 145
2 1 4 0 0 0 12 15 17 0 0 2
87 66
65 66
2 1 4 0 0 8320 12 19 17 0 0 3
85 103
65 103
65 66
1 2 2 0 0 0 0 10 11 0 0 2
328 87
328 86
1 2 2 0 0 0 0 13 12 0 0 2
328 133
328 132
2 1 2 0 0 4224 0 17 16 0 0 2
23 66
13 66
1 3 2 0 0 0 0 14 15 0 0 2
87 75
87 74
1 3 2 0 0 0 0 18 19 0 0 2
85 112
85 111
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
