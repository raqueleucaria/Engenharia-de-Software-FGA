CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 30 400 10
176 80 1918 940
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
47 C:\Users\User\Desktop\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
20
7 Ground~
168 327 148 0 1 3
0 9
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9424 0 0
2
44773.7 0
0
4 LED~
171 327 132 0 2 2
10 3 9
0
0 0 864 0
4 LED0
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
9968 0 0
2
44773.7 0
0
9 Inverter~
13 136 177 0 2 22
0 7 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
9281 0 0
2
44773.7 0
0
9 Inverter~
13 135 143 0 2 22
0 9 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
8464 0 0
2
44773.7 0
0
9 Inverter~
13 134 107 0 2 22
0 9 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
7168 0 0
2
44773.7 0
0
9 Inverter~
13 136 70 0 2 22
0 9 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3171 0 0
2
44773.7 0
0
8 3-In OR~
219 279 122 0 4 22
0 13 14 12 3
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
4139 0 0
2
44773.7 0
0
5 7415~
219 206 164 0 4 22
0 10 5 4 12
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 1 0
1 U
6435 0 0
2
44773.7 0
0
5 7415~
219 206 122 0 4 22
0 10 6 5 14
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
5283 0 0
2
44773.7 0
0
5 7415~
219 206 79 0 4 22
0 10 6 4 13
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 1 0
1 U
6874 0 0
2
44773.7 0
0
7 Ground~
168 87 81 0 1 3
0 9
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5305 0 0
2
44773.7 1
0
12 SPDT Switch~
164 104 70 0 3 11
0 9 7 9
0
0 0 4720 0
0
1 M
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
34 0 0
2
44773.7 0
0
7 Ground~
168 87 188 0 1 3
0 9
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
969 0 0
2
44773.7 1
0
12 SPDT Switch~
164 104 177 0 10 11
0 7 7 9 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 F3
-7 -16 7 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
8402 0 0
2
44773.7 0
0
7 Ground~
168 87 154 0 1 3
0 9
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3751 0 0
2
44773.7 1
0
12 SPDT Switch~
164 104 143 0 3 11
0 9 7 9
0
0 0 4720 0
0
2 F2
-7 -16 7 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
4292 0 0
2
44773.7 0
0
7 Ground~
168 13 72 0 1 3
0 9
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6118 0 0
2
5.90041e-315 0
0
9 V Source~
197 45 65 0 2 5
0 7 9
0
0 0 17264 270
2 5V
-7 -20 7 -12
3 Vs1
-11 -30 10 -22
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
34 0 0
2
5.90041e-315 0
0
7 Ground~
168 85 118 0 1 3
0 9
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6357 0 0
2
5.90041e-315 0
0
12 SPDT Switch~
164 102 107 0 3 11
0 9 7 9
0
0 0 4720 0
0
2 F1
-7 -16 7 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
319 0 0
2
5.90041e-315 0
0
27
1 2 9 0 0 0 2 1 2 0 0 2
327 142
327 142
4 1 3 0 0 4224 0 7 2 0 0 2
312 122
327 122
3 0 4 0 0 4096 0 8 0 0 7 2
182 173
162 173
0 2 5 0 0 4224 0 0 8 5 0 3
155 131
155 164
182 164
2 3 5 0 0 0 0 5 9 0 0 3
155 107
155 131
182 131
2 0 6 0 0 4096 0 9 0 0 8 2
182 122
166 122
3 2 4 0 0 8320 0 10 3 0 0 4
182 88
162 88
162 177
157 177
2 2 6 0 0 8320 0 4 10 0 0 4
156 143
166 143
166 79
182 79
1 1 7 0 0 0 0 3 14 0 0 2
121 177
121 177
1 1 9 0 0 4224 8 4 16 0 0 2
120 143
121 143
1 1 9 0 0 0 0 5 20 0 0 2
119 107
119 107
2 0 10 0 0 8320 0 6 0 0 13 3
157 70
172 70
172 114
1 1 10 0 0 0 0 8 9 0 0 4
182 155
172 155
172 113
182 113
2 1 10 0 0 0 0 6 10 0 0 2
157 70
182 70
1 1 9 0 0 0 11 6 12 0 0 2
121 70
121 70
4 3 12 0 0 8320 0 8 7 0 0 3
227 164
227 131
266 131
4 1 13 0 0 8320 0 10 7 0 0 3
227 79
227 113
266 113
4 2 14 0 0 4224 0 9 7 0 0 2
227 122
267 122
2 0 7 0 0 4096 15 12 0 0 22 2
87 66
65 66
2 0 7 0 0 0 15 20 0 0 22 2
85 103
65 103
2 0 7 0 0 0 15 16 0 0 22 2
87 139
65 139
1 2 7 0 0 4224 15 18 14 0 0 3
65 66
65 173
87 173
2 1 9 0 0 4224 2 18 17 0 0 2
23 66
13 66
1 3 9 0 0 0 2 11 12 0 0 2
87 75
87 74
1 3 9 0 0 0 2 13 14 0 0 2
87 182
87 181
1 3 9 0 0 0 2 15 16 0 0 2
87 148
87 147
1 3 9 0 0 0 2 19 20 0 0 2
85 112
85 111
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
