CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 70 30 400 10
176 80 1918 940
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
47 C:\Users\User\Desktop\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
8 2-In OR~
219 200 117 0 3 22
0 3 4 8
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3472 0 0
2
44774.5 0
0
9 3-In AND~
219 148 174 0 4 22
0 7 7 7 4
0
0 0 624 0
5 74F11
-18 -28 17 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 1 0
1 U
9998 0 0
2
44774.5 0
0
12 SPDT Switch~
164 103 259 0 10 11
0 7 7 3 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 D
-4 -15 3 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
3536 0 0
2
44774.4 1
0
7 Ground~
168 86 269 0 1 3
0 3
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
44774.4 0
0
7 Ground~
168 32 188 0 1 3
0 3
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3835 0 0
2
44774.4 0
0
9 V Source~
197 32 162 0 2 5
0 7 3
0
0 0 17264 0
2 5V
16 0 30 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
3670 0 0
2
44774.4 1
0
7 Ground~
168 234 194 0 1 3
0 3
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5616 0 0
2
44774.4 2
0
7 Ground~
168 84 227 0 1 3
0 3
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9323 0 0
2
44774.4 3
0
7 Ground~
168 84 175 0 1 3
0 3
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
317 0 0
2
44774.4 4
0
7 Ground~
168 85 118 0 1 3
0 3
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3108 0 0
2
44774.4 5
0
12 SPDT Switch~
164 101 217 0 10 11
0 7 7 3 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 C
-4 -15 3 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
4299 0 0
2
44774.4 6
0
12 SPDT Switch~
164 101 165 0 10 11
0 7 7 3 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 B
-4 -15 3 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9672 0 0
2
44774.4 7
0
12 SPDT Switch~
164 102 108 0 3 11
0 3 7 3
0
0 0 4720 0
0
1 A
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
7876 0 0
2
44774.4 8
0
4 LED~
171 234 178 0 2 2
10 8 3
0
0 0 496 0
4 LED1
13 0 41 8
0
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6369 0 0
2
44774.4 9
0
16
1 1 3 0 0 4224 0 13 1 0 0 2
119 108
187 108
2 4 4 0 0 8320 0 1 2 0 0 3
187 126
169 126
169 174
3 1 7 0 0 4224 5 2 3 0 0 3
124 183
124 259
120 259
2 1 7 0 0 8320 6 2 11 0 0 3
124 174
118 174
118 217
1 1 7 0 0 4224 0 2 12 0 0 2
124 165
118 165
3 1 8 0 0 8336 0 1 14 0 0 3
233 117
234 117
234 168
2 0 7 0 0 4096 9 11 0 0 9 2
84 213
67 213
2 0 7 0 0 0 9 12 0 0 9 2
84 161
67 161
2 0 7 0 0 8320 9 3 0 0 12 3
86 255
67 255
67 104
1 3 3 0 0 0 2 4 3 0 0 2
86 263
86 263
1 2 3 0 0 0 2 7 14 0 0 2
234 188
234 188
2 1 7 0 0 128 9 13 6 0 0 3
85 104
32 104
32 141
1 2 3 0 0 4224 2 5 6 0 0 2
32 182
32 183
1 3 3 0 0 0 2 8 11 0 0 2
84 221
84 221
1 3 3 0 0 0 2 9 12 0 0 2
84 169
84 169
1 3 3 0 0 0 2 10 13 0 0 2
85 112
85 112
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
