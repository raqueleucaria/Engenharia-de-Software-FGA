CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 60 30 200 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
47 C:\Users\User\Desktop\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
44
7 Ground~
168 464 416 0 1 3
0 2
0
0 0 53344 90
0
5 GND14
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5130 0 0
2
44777 0
0
7 Ground~
168 454 287 0 1 3
0 2
0
0 0 53344 90
0
5 GND13
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
391 0 0
2
44777 0
0
4 LED~
171 444 416 0 1 2
10 11
0
0 0 880 90
4 LED0
-12 -21 16 -13
2 U7
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3124 0 0
2
44777 0
0
4 LED~
171 434 287 0 1 2
10 11
0
0 0 880 90
4 LED0
-12 -21 16 -13
2 U6
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3421 0 0
2
44777 0
0
9 Inverter~
13 250 505 0 2 22
0 5 15
0
0 0 96 0
6 74LS04
-21 -19 21 -11
2 AF
-7 -29 7 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 512 6 6 6 0
1 U
8157 0 0
2
44777 0
0
9 Inverter~
13 243 395 0 2 22
0 5 15
0
0 0 96 0
6 74LS04
-21 -19 21 -11
2 AE
-7 -29 7 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 512 6 5 6 0
1 U
5572 0 0
2
44777 0
0
9 Inverter~
13 244 335 0 2 22
0 5 15
0
0 0 96 0
6 74LS04
-21 -19 21 -11
2 AD
-7 -29 7 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 512 6 4 6 0
1 U
8901 0 0
2
44777 0
0
7 Ground~
168 44 405 0 1 3
0 2
0
0 0 53344 0
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7361 0 0
2
44776.9 0
0
7 Ground~
168 110 480 0 1 3
0 2
0
0 0 53344 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4747 0 0
2
44776.9 0
0
7 Ground~
168 111 404 0 1 3
0 2
0
0 0 53344 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
972 0 0
2
44776.9 0
0
7 Ground~
168 108 345 0 1 3
0 2
0
0 0 53344 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3472 0 0
2
44776.9 0
0
7 Ground~
168 108 286 0 1 3
0 2
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9998 0 0
2
44776.9 0
0
8 3-In OR~
219 405 417 0 1 22
0 0
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U2B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 7 0
1 U
3536 0 0
2
44776.9 0
0
5 4073~
219 304 496 0 1 22
0 0
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 9 0
1 U
4597 0 0
2
44776.9 0
0
5 4073~
219 306 415 0 1 22
0 0
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 9 0
1 U
3835 0 0
2
44776.9 0
0
5 4073~
219 306 345 0 1 22
0 0
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 9 0
1 U
3670 0 0
2
44776.9 0
0
5 4012~
219 400 288 0 1 22
0 0
0
0 0 608 0
4 4012
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 8 0
1 U
5616 0 0
2
44776.9 0
0
12 SPDT Switch~
164 126 470 0 1 11
0 0
0
0 0 4704 0
0
2 S4
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
9323 0 0
2
44776.9 0
0
12 SPDT Switch~
164 127 395 0 1 11
0 0
0
0 0 4704 0
0
2 S3
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
317 0 0
2
44776.9 0
0
12 SPDT Switch~
164 124 335 0 1 11
0 0
0
0 0 4704 0
0
2 S2
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
3108 0 0
2
44776.9 0
0
12 SPDT Switch~
164 124 276 0 1 11
0 0
0
0 0 4704 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
4299 0 0
2
44776.9 0
0
9 V Source~
197 44 379 0 1 5
0 0
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs2
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
9672 0 0
2
44776.9 0
0
8 3-In OR~
219 287 163 0 4 22
0 10 9 8 7
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 7 0
1 U
7876 0 0
2
5.90041e-315 0
0
9 Inverter~
13 201 196 0 2 22
0 5 13
0
0 0 112 0
6 74LS04
-21 -19 21 -11
2 A1
-7 -29 7 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 3 6 0
1 U
6369 0 0
2
5.90041e-315 0
0
9 Inverter~
13 201 154 0 2 22
0 5 14
0
0 0 112 0
6 74LS04
-21 -19 21 -11
2 A2
-7 -29 7 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 2 6 0
1 U
9172 0 0
2
5.90041e-315 0
0
9 Inverter~
13 201 113 0 2 22
0 5 15
0
0 0 112 0
6 74LS04
-21 -19 21 -11
2 A3
-7 -29 7 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 90
65 0 0 512 6 1 6 0
1 U
7100 0 0
2
5.90041e-315 0
0
5 7415~
219 244 205 0 4 22
0 16 5 5 8
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 512 3 3 5 0
1 U
3820 0 0
2
5.90041e-315 0
0
5 7415~
219 244 163 0 4 22
0 17 5 5 9
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 512 3 2 5 0
1 U
7678 0 0
2
5.90041e-315 0
0
5 7415~
219 244 122 0 4 22
0 18 5 5 10
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 512 3 1 5 0
1 U
961 0 0
2
5.90041e-315 0
0
4 LED~
171 329 182 0 2 2
10 7 2
0
0 0 880 0
4 LED0
17 0 45 8
1 M
27 -10 34 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3178 0 0
2
5.90041e-315 5.26354e-315
0
7 Ground~
168 329 198 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3409 0 0
2
5.90041e-315 0
0
9 4-In AND~
219 305 83 0 5 22
0 5 5 5 5 11
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U4A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 4 0
1 U
3951 0 0
2
5.90041e-315 0
0
7 Ground~
168 327 123 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8885 0 0
2
5.90041e-315 0
0
4 LED~
171 327 108 0 2 2
10 11 2
0
0 0 880 0
4 LED0
17 0 45 8
1 U
28 -10 35 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3780 0 0
2
5.90041e-315 0
0
7 Ground~
168 87 81 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9265 0 0
2
5.90041e-315 5.26354e-315
0
12 SPDT Switch~
164 104 70 0 10 11
0 5 5 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 A
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9442 0 0
2
5.90041e-315 0
0
7 Ground~
168 87 188 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9424 0 0
2
5.90041e-315 5.26354e-315
0
12 SPDT Switch~
164 104 177 0 10 11
0 5 5 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 D
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9968 0 0
2
5.90041e-315 0
0
7 Ground~
168 87 154 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9281 0 0
2
5.90041e-315 5.26354e-315
0
12 SPDT Switch~
164 104 143 0 10 11
0 5 5 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 C
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
8464 0 0
2
5.90041e-315 0
0
7 Ground~
168 13 72 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7168 0 0
2
44776.9 0
0
9 V Source~
197 45 65 0 2 5
0 5 2
0
0 0 17264 270
2 5V
-7 -20 7 -12
3 Vs1
-11 -30 10 -22
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
3171 0 0
2
44776.9 1
0
7 Ground~
168 85 118 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4139 0 0
2
44776.9 2
0
12 SPDT Switch~
164 102 107 0 10 11
0 5 5 2 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 B
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
6435 0 0
2
44776.9 3
0
64
1 2 0 0 0 0 0 1 3 0 0 2
457 417
457 417
2 1 0 0 0 0 0 4 2 0 0 2
447 288
447 288
4 1 0 0 0 0 0 13 3 0 0 2
438 417
437 417
5 1 0 0 0 0 0 17 4 0 0 2
427 288
427 288
4 3 0 0 0 0 0 14 13 0 0 4
325 496
354 496
354 426
392 426
4 1 0 0 0 0 0 16 13 0 0 4
327 345
354 345
354 408
392 408
2 4 0 0 0 0 0 13 15 0 0 3
393 417
393 415
327 415
2 3 0 0 0 0 0 5 14 0 0 2
271 505
280 505
2 1 0 0 0 0 0 6 15 0 0 3
264 395
282 395
282 406
2 1 0 0 0 0 0 7 16 0 0 3
265 335
282 335
282 336
3 0 0 0 0 0 0 16 0 0 16 2
282 354
199 354
0 1 0 0 0 0 0 0 5 16 0 3
199 470
199 505
235 505
0 1 0 0 0 0 0 0 14 14 0 3
180 395
180 487
280 487
0 1 0 0 0 0 0 0 6 15 0 2
179 395
228 395
1 3 0 0 0 0 0 19 17 0 0 4
144 395
179 395
179 293
376 293
1 4 0 0 0 0 0 18 17 0 0 4
143 470
199 470
199 302
376 302
3 0 0 0 0 0 0 15 0 0 18 3
282 424
157 424
157 335
1 1 0 0 0 0 0 20 7 0 0 2
141 335
229 335
1 2 0 0 0 0 0 20 17 0 0 4
141 335
157 335
157 284
376 284
2 0 0 0 0 0 0 15 0 0 22 4
282 415
220 415
220 414
205 414
2 0 0 0 0 0 0 16 0 0 22 2
282 345
205 345
0 2 0 0 0 0 0 0 14 23 0 3
205 274
205 496
280 496
1 1 0 0 0 0 0 21 17 0 0 5
141 276
141 274
205 274
205 275
376 275
0 2 0 0 0 0 0 0 18 25 0 3
86 390
86 466
109 466
0 2 0 0 0 0 0 0 19 26 0 3
86 330
86 391
110 391
0 2 0 0 0 0 0 0 20 27 0 3
86 272
86 331
107 331
1 2 0 0 0 0 0 22 21 0 0 3
44 358
44 272
107 272
1 2 0 0 0 0 0 8 22 0 0 2
44 399
44 400
1 3 0 0 0 0 0 9 18 0 0 2
110 474
109 474
1 3 0 0 0 0 0 10 19 0 0 3
111 398
111 399
110 399
1 3 0 0 0 0 0 11 20 0 0 2
108 339
107 339
1 3 0 0 0 0 0 12 21 0 0 2
108 280
107 280
2 1 0 0 0 0 0 26 29 0 0 2
222 113
220 113
2 1 0 0 0 0 0 25 28 0 0 2
222 154
220 154
2 1 0 0 0 0 0 24 27 0 0 2
222 196
220 196
3 0 5 0 0 8192 3 27 0 0 48 3
220 214
170 214
170 154
0 2 5 0 0 8192 4 0 27 39 0 3
157 163
157 205
220 205
3 0 5 0 0 4096 0 28 0 0 49 3
220 172
142 172
142 113
0 2 5 0 0 0 4 0 28 41 0 3
157 122
157 163
220 163
3 0 5 0 0 4096 6 29 0 0 50 3
220 131
148 131
148 97
2 0 5 0 0 4096 4 29 0 0 53 3
220 122
156 122
156 70
1 2 2 0 0 4096 0 33 34 0 0 2
327 117
327 118
4 1 7 0 0 4224 0 23 30 0 0 3
320 163
329 163
329 172
4 3 8 0 0 8320 0 27 23 0 0 3
265 205
274 205
274 172
4 2 9 0 0 4224 0 28 23 0 0 2
265 163
275 163
4 1 10 0 0 8320 0 29 23 0 0 3
265 122
274 122
274 154
1 1 5 0 0 0 6 24 38 0 0 3
186 196
121 196
121 177
1 1 5 0 0 4096 3 25 40 0 0 3
186 154
121 154
121 143
1 1 5 0 0 0 0 44 26 0 0 3
119 107
119 113
186 113
1 4 5 0 0 12416 6 38 32 0 0 4
121 177
132 177
132 97
281 97
1 3 5 0 0 12416 3 40 32 0 0 4
121 143
126 143
126 88
281 88
1 2 5 0 0 8320 0 44 32 0 0 3
119 107
119 79
281 79
1 1 5 0 0 4224 4 36 32 0 0 2
121 70
281 70
5 1 11 0 0 8320 0 32 34 0 0 3
326 83
327 83
327 98
1 2 2 0 0 0 0 31 30 0 0 2
329 192
329 192
2 0 5 0 0 4096 12 36 0 0 59 2
87 66
65 66
2 0 5 0 0 0 12 44 0 0 59 2
85 103
65 103
2 0 5 0 0 0 12 40 0 0 59 2
87 139
65 139
1 2 5 0 0 4224 12 42 38 0 0 3
65 66
65 173
87 173
2 1 2 0 0 4224 0 42 41 0 0 2
23 66
13 66
1 3 2 0 0 0 0 35 36 0 0 2
87 75
87 74
1 3 2 0 0 0 0 37 38 0 0 2
87 182
87 181
1 3 2 0 0 0 0 39 40 0 0 2
87 148
87 147
1 3 2 0 0 0 0 43 44 0 0 2
85 112
85 111
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
