CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 400 10
176 80 1918 940
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
47 C:\Users\User\Desktop\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
13
9 Inverter~
13 165 121 0 2 22
0 3 6
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
8402 0 0
2
44774.4 0
0
9 Inverter~
13 165 88 0 2 22
0 7 8
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3751 0 0
2
44774.4 0
0
9 2-In AND~
219 210 79 0 3 22
0 3 8 5
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4292 0 0
2
44774.4 0
0
7 Ground~
168 328 93 0 1 3
0 7
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6118 0 0
2
44773.8 1
0
4 LED~
171 328 76 0 2 2
10 5 7
0
0 0 864 0
4 LED0
22 22 50 30
2 VE
25 -10 39 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
34 0 0
2
44773.8 0
0
4 LED~
171 328 122 0 2 2
10 6 7
0
0 0 864 0
4 LED0
22 22 50 30
2 VS
25 -10 39 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6357 0 0
2
5.90041e-315 0
0
7 Ground~
168 328 139 0 1 3
0 7
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
319 0 0
2
5.90041e-315 0
0
7 Ground~
168 87 81 0 1 3
0 7
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3976 0 0
2
5.90041e-315 5.26354e-315
0
12 SPDT Switch~
164 104 70 0 10 11
0 3 3 7 0 0 0 0 0 0
1
0
0 0 4720 0
0
1 I
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
7634 0 0
2
5.90041e-315 0
0
7 Ground~
168 13 72 0 1 3
0 7
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
523 0 0
2
44773.8 0
0
9 V Source~
197 45 65 0 2 5
0 3 7
0
0 0 17264 270
2 5V
-7 -20 7 -12
3 Vs1
-11 -30 10 -22
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
6748 0 0
2
44773.8 1
0
7 Ground~
168 85 118 0 1 3
0 7
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6901 0 0
2
44773.8 2
0
12 SPDT Switch~
164 102 107 0 3 11
0 7 3 7
0
0 0 4720 0
0
1 A
-4 -16 3 -8
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
842 0 0
2
44773.8 3
0
13
1 0 3 0 0 8192 0 1 0 0 3 3
150 121
131 121
131 70
2 1 3 0 0 4096 4 9 11 0 0 2
87 66
65 66
1 1 3 0 0 4224 0 9 3 0 0 2
121 70
186 70
3 1 5 0 0 4224 0 3 5 0 0 4
231 79
311 79
311 66
328 66
1 2 6 0 0 4224 0 6 1 0 0 3
328 112
186 112
186 121
1 1 7 0 0 4224 0 13 2 0 0 3
119 107
150 107
150 88
2 2 8 0 0 0 0 2 3 0 0 2
186 88
186 88
2 1 3 0 0 8320 4 13 11 0 0 3
85 103
65 103
65 66
1 2 7 0 0 4112 2 4 5 0 0 2
328 87
328 86
1 2 7 0 0 0 2 7 6 0 0 2
328 133
328 132
2 1 7 0 0 4224 2 11 10 0 0 2
23 66
13 66
1 3 7 0 0 0 2 8 9 0 0 2
87 75
87 74
1 3 7 0 0 0 2 12 13 0 0 2
85 112
85 111
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
